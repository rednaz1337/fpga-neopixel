module rainbow();

endmodule